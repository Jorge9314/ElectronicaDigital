library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity motores is
    Port ( CLK : in  STD_LOGIC;
           Salida : out  STD_LOGIC_VECTOR (0 downto 3);
           Entrada : in  STD_LOGIC);
end motores;

architecture Behavioral of motores is

begin


end Behavioral;

